-- Library & Use Statements
-- Entity Declaration 

-- Architecture Declaration�
�   -- Component Declaration 
    -- Signals & Constants Declaration�
-- Begin Architecture

    -------------------------------------------
    -- Instantiation DUT (Device under Test)
    -------------------------------------------
	-- Clock Generation Process (with wait)
    -------------------------------------------
    -- Stimuli and Check Process (with wait & ASSERT)
	-------------------------------------------

�-- End Architecture 
