-- Library & Use Statements
-- Entity Declaration 

-- Architecture Declaration�
�   -- Components Declaration 
    -- Signals & Constants Declaration
	�
-- Begin Architecture

    -------------------------------------------
    -- Instantiation Block - 1
    -------------------------------------------
	-- Instantiation Block � 2 ...
    -------------------------------------------
    -- Concurrent Assignments  
    -- e.g. Assign outputs from intermediate signals
	-------------------------------------------

�-- End Architecture 
