-------------------------------------------------------------------------------
--  _____       ______  _____                                                 -
-- |_   _|     |  ____|/ ____|                                                -
--   | |  _ __ | |__  | (___    Institute of Embedded Systems                 -
--   | | | '_ \|  __|  \___ \   Zuercher Hochschule Winterthur                -
--  _| |_| | | | |____ ____) |  (University of Applied Sciences)              -
-- |_____|_| |_|______|_____/   8401 Winterthur, Switzerland                  -             
-------------------------------------------------------------------------------
--
-- Project     : HDMI_TEA
-- Description : debounce.vhd
--
-- $LastChangedDate$
-- $Rev$
-- $Author$
-------------------------------------------------------------------------------
-- Change History
-- Date     |Name      |Modification
------------|----------|-------------------------------------------------------
-- 21.05.15 | scln     | file created
-- 05.06.15 | scln     | changed reset values to '1'
-------------------------------------------------------------------------------


-------------------------------------------------------------------------------
-- Package / Component Declaration
-------------------------------------------------------------------------------
-- Include in Design:
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

-------------------------------------------------------------------------------
-- Architecture
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;


entity debounce is
		PORT(
			clk_100M		: IN    std_logic;
			reset_n			: IN    std_logic;
			signal_in		: IN    std_logic;
			signal_out		: OUT   std_logic
		);
end entity;


-- begin of Architecture
architecture rtl of debounce is

-------------------------------------------------------------------------------
-- Constant declaration
-------------------------------------------------------------------------------


---------------------------------------------------------------------------------
---- Components
---------------------------------------------------------------------------------


---------------------------------------------------------------------------------
---- Signal declaration
---------------------------------------------------------------------------------
SIGNAL Q1, Q2, Q3	: std_logic := '1';

BEGIN
---------------------------------------------------------------------------------
---- Components initiation
---------------------------------------------------------------------------------
gen_clk: PROCESS (clk_100M, reset_n)
BEGIN
	
	IF reset_n = '0' THEN
		Q1 <= '1';
		Q2 <= '1';
		Q3 <= '1';
	ELSIF rising_edge(clk_100M) THEN
		Q1 <= signal_in;
		Q2 <= Q1;
		Q3 <= Q2;
	END IF;

END PROCESS gen_clk;
---------------------------------------------------------------------------------
---- Signal initiation                                          
---------------------------------------------------------------------------------

signal_out <= Q1 AND Q2 AND Q3;
	
end architecture;

