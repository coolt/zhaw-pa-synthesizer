-- Library & Use Statements

-- Entity Declaration 

-- Architecture Declaration�
-- Signals & Constants Declaration�
-- Begin Architecture

    -------------------------------------------
    -- Process for combinatorial logic
    -------------------------------------------
	-- Process for registers (flip-flops)
    -------------------------------------------
    -- Concurrent Assignements  
    -- e.g. Assign outputs from intermediate signals
	-------------------------------------------

�-- End Architecture 
